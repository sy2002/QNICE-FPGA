----------------------------------------------------------------------------------
-- EAE - Extended Arithmetic Element inspired by the PDP-11
-- 
-- done in May 2016 by sy2002
----------------------------------------------------------------------------------

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity EAE is
end EAE;

architecture Behavioral of EAE is

begin


end Behavioral;

